//-------------------------------------------------------------------------
//						www.verificationguide.com
//-------------------------------------------------------------------------
interface intf(input logic clk,reset);
  
  //declaring the signals
  logic [1:0] opcode;
  logic [3:0] a;
  logic [3:0] b;
  logic [8:0] c;
  
endinterface
